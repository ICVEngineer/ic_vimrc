Vim�UnDo� ����p�mR����ol0r�H���)	�gH2�   -                                      W��    _�                             ����                                                                                                                                                                                                                                                                                                                                                             W��     �                  lab5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             W��     �                   5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             W��0     �                module hello_world();5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             W��7     �               begin5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             W��;     �               begin5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             W��D     �                   $display();5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             W��F    �                   $display("");5�_�                           ����                                                                                                                                                                                                                                                                                                                                                             W��R    �                   $display("hello world!");5�_�         
             	    ����                                                                                                                                                                                                                                                                                                                                                 v       W���    �                  �               �                 	endmodule5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       W���     �                   �             �             5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       W���     �                �             �             5�_�                           ����                                                                                                                                                                                                                                                                                                                                                v       W���    �                �             �             5�_�                           ����                                                                                                                                                                                                                                                                                                                                         $       v   $    W���    �                �             �             5�_�                      9    ����                                                                                                                                                                                                                                                                                                                                                         W�
�   	 �      	         9 that is used more often on MS-Windows than on X-Windows.5�_�                           ����                                                                                                                                                                                                                                                                                                                                                         W�    
 �      	         > that is used more often on MS-Windows than on X-Windows.     5�_�                       $    ����                                                                                                                                                                                                                                                                                                                            	          	                 W��     �               $Visual mode, because it is also used5�_�                             ����                                                                                                                                                                                                                                                                                                                            	          	                 W��     �             �             5�_�                              ����                                                                                                                                                                                                                                                                                                                                         2          2    W��    �                  �               5�_�                     L    ����                                                                                                                                                                                                                                                                                                                                                         W�
�     �             �               ^But both can do it.  You already know about Visual mode.  Select mode is likee often on MS-Win   ^Visual mode, because it is also used to select text.  But there is an obviousit.  You already    ^difference: When typi                                                        ause it is also u   R is used more often on MS-Windows than on X-Windows.                          typi   ^But both can do it.  You already know about Visual mode.  Select mode is liketen on MS-Windows   MVisual mode, because it is also used to select text.  But there is an obvious5�_�                        ]    ����                                                                                                                                                                                                                                                                                                                                                         W�
�     �             �               oBut both can do it.  You already know about Visual mode.  Select mode is likee often on MS-Wine often on MS-Win   oVisual mode, because it is also used to select text.  But there is an obviousit.  You already it.  You already    odifference: When typi                                                        ause it is also uause it is also u   c is used more often on MS-Windows than on X-Windows.                          typi             typi   oBut both can do it.  You already know about Visual mode.  Select mode is liketen on MS-Windowsten on MS-Windows   MVisual mode, because it is also used to select text.  But there is an obvious5�_�                      L    ����                                                                                                                                                                                                                                                                                                                                                         W�
�     �             �               ^But both can do it.  You already know about Visual mode.  Select mode is likee often on MS-Win   ^Visual mode, because it is also used to select text.  But there is an obviousit.  You already    ^difference: When typi                                                        ause it is also u   R is used more often on MS-Windows than on X-Windows.                          typi   ^But both can do it.  You already know about Visual mode.  Select mode is liketen on MS-Windows   MVisual mode, because it is also used to select text.  But there is an obvious5�_�                      L    ����                                                                                                                                                                                                                                                                                                                                                         W�
�     �             �               ^But both can do it.  You already know about Visual mode.  Select mode is likee often on MS-Win   ^Visual mode, because it is also used to select text.  But there is an obviousit.  You already    ^difference: When typi                                                        ause it is also u   R is used more often on MS-Windows than on X-Windows.                          typi   ^But both can do it.  You already know about Visual mode.  Select mode is liketen on MS-Windows   MVisual mode, because it is also used to select text.  But there is an obvious5�_�                     L    ����                                                                                                                                                                                                                                                                                                                                                         W�
�     �             �               ^But both can do it.  You already know about Visual mode.  Select mode is likee often on MS-Win   ^Visual mode, because it is also used to select text.  But there is an obviousit.  You already    ^difference: When typi                                                        ause it is also u   R is used more often on MS-Windows than on X-Windows.                          typi   ^But both can do it.  You already know about Visual mode.  Select mode is liketen on MS-Windows   MVisual mode, because it is also used to select text.  But there is an obvious5�_�                        M    ����                                                                                                                                                                                                                                                                                                                                                         W�
�     �             �               oBut both can do it.  You already know about Visual mode.  Select mode is likeee often on MS-Win often on MS-Win   oVisual mode, because it is also used to select text.  But there is an obviousiit.  You already t.  You already    odifference: When typi                                                        aause it is also uuse it is also u   c is used more often on MS-Windows than on X-Windows.                           typi            typi   oBut both can do it.  You already know about Visual mode.  Select mode is liketten on MS-Windowsen on MS-Windows   MVisual mode, because it is also used to select text.  But there is an obvious5�_�                      7    ����                                                                                                                                                                                                                                                                                                                                                         W�
�     �             �               I     is used more often on MS-Windows than on X-Windows.e often on MS-Win   ^But both can do it.  You already know about Visual mode.it.  You already   Select mode is like   ^Visual mode, because it is also used to select text.  Buause it is also ut there is an obvious   =difference: When typi                                    typi   I is used more often on MS-Windows than on X-Windows.    ten on MS-Windows   MBut both can do it.  You already know about Visual mode.  Select mode is like5�_�                   	   &    ����                                                                                                                                                                                                                                                                                                                                                             W�
j     �      	          5�_�                   	   &    ����                                                                                                                                                                                                                                                                                                                                                             W�
g     �   	   
          5�_�                          ����                                                                                                                                                                                                                                                                                                                                                             W�
^     �              5�_�                             ����                                                                                                                                                                                                                                                                                                                                                             W�
_     �              5�_�         	      
          ����                                                                                                                                                                                                                                                                                                                                                 v       W���     �                   $pisplay("hello world!");5�_�   
                         ����                                                                                                                                                                                                                                                                                                                                                 v       W���     �             �                   $pdisplay("hello world!");5�_�              
   	           ����                                                                                                                                                                                                                                                                                                                                                             W��:     �                initiel�                    $displey("hello world!");5��